module transmitter (
   
);
  
endmodule
